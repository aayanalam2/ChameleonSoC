module or2 (
    input wire A, B,  // Inputs
    output wire Y     // Output
);
    assign Y = A | B; // OR operation
endmodule

